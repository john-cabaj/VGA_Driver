library verilog;
use verilog.vl_types.all;
entity t_timing_generator is
end t_timing_generator;
