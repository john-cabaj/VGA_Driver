library verilog;
use verilog.vl_types.all;
entity t_display_plane is
end t_display_plane;
